//`define define  
// 4.3' 480*272
`define  H_SYNC_4342     11'd41
`define  H_BACK_4342     11'd2
`define  H_DISP_4342     11'd480    
`define  H_FRONT_4342    11'd2
`define  H_TOTAL_4342    11'd525
   
`define  V_SYNC_4342     11'd10     
`define  V_BACK_4342     11'd2      
`define  V_DISP_4342     11'd272    
`define  V_FRONT_4342    11'd2      
`define  V_TOTAL_4342    11'd286
   
// 7' 800*480   
`define  H_SYNC_7084     11'd128
`define  H_BACK_7084     11'd88
`define  H_DISP_7084     11'd800
`define  H_FRONT_7084    11'd40
`define  H_TOTAL_7084    11'd1056
   
`define  V_SYNC_7084     11'd2
`define  V_BACK_7084     11'd33
`define  V_DISP_7084     11'd480
`define  V_FRONT_7084    11'd10
`define  V_TOTAL_7084    11'd525
   
// 7' 1024*600   
`define  H_SYNC_7016     11'd20
`define  H_BACK_7016     11'd140
`define  H_DISP_7016     11'd1024
`define  H_FRONT_7016    11'd160
`define  H_TOTAL_7016    11'd1344
   
`define  V_SYNC_7016     11'd3
`define  V_BACK_7016     11'd20
`define  V_DISP_7016     11'd600
`define  V_FRONT_7016    11'd12
`define  V_TOTAL_7016    11'd635
   
// 10.1' 1280*800   
`define  H_SYNC_1018     11'd10
`define  H_BACK_1018     11'd80
`define  H_DISP_1018     11'd1280
`define  H_FRONT_1018    11'd70
`define  H_TOTAL_1018    11'd1440
   
`define  V_SYNC_1018     11'd3
`define  V_BACK_1018     11'd10
`define  V_DISP_1018     11'd800
`define  V_FRONT_1018    11'd10
`define  V_TOTAL_1018    11'd823

// 4.3' 800*480   
`define  H_SYNC_4384     11'd128
`define  H_BACK_4384     11'd88
`define  H_DISP_4384     11'd800
`define  H_FRONT_4384    11'd40
`define  H_TOTAL_4384    11'd1056
   
`define  V_SYNC_4384     11'd2
`define  V_BACK_4384     11'd33
`define  V_DISP_4384     11'd480
`define  V_FRONT_4384    11'd10
`define  V_TOTAL_4384    11'd525